// PyXHDL support functions.
