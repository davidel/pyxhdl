/* verilator lint_off WIDTH */

`timescale @{TS_INT:1} @{TIME_UNIT:ns} / @{TS_RES:1} ps
