/* verilator lint_off WIDTH */

`timescale 1 ns / 100 ps


package fp;
  let MAX(A, B) = ((A > B) ? A : B);
  let MIN(A, B) = ((A > B) ? B : A);
  let ABS(A) = (($signed(A) >= 0) ? A : -$signed(A));
  let FABS(A) = ((A >= 0.0) ? A : -A);

  let EXP_OFFSET(NX) = (2**(NX - 1) - 1);
endpackage

// This in theory should be a typedef within the FPU interface, but then
// many HDL tools do not support hierarchical type dereferencing.
`define IEEE754(NX, NM) \
struct packed { \
  logic  sign; \
  logic [NX - 1: 0] exp; \
  logic [NM - 1: 0] mant; \
  }


// PyXHDL support functions.

// Entity "MatMult" is "MatMult" with:
// 	args={'A': 'uint(4, 4, 16)', 'B': 'uint(4, 4, 16)', 'XOUT': 'uint(4, 4, 16)'}
// 	kwargs={}
module MatMult(A, B, XOUT);
  input logic [15: 0] A[4][4];
  input logic [15: 0] B[4][4];
  output logic [15: 0] XOUT[4][4];
  logic [15: 0] XOUT_[4][4];
  always @(A or B)
  mat_mult : begin
    XOUT_[0][0] = (((0 + 16'(A[0][0] * B[0][0])) + 16'(A[0][1] * B[1][0])) + 16'(A[0][2] * B[2][0])) + 16'(A[0][3] * B[3][0]);
    XOUT_[0][1] = (((0 + 16'(A[0][0] * B[0][1])) + 16'(A[0][1] * B[1][1])) + 16'(A[0][2] * B[2][1])) + 16'(A[0][3] * B[3][1]);
    XOUT_[0][2] = (((0 + 16'(A[0][0] * B[0][2])) + 16'(A[0][1] * B[1][2])) + 16'(A[0][2] * B[2][2])) + 16'(A[0][3] * B[3][2]);
    XOUT_[0][3] = (((0 + 16'(A[0][0] * B[0][3])) + 16'(A[0][1] * B[1][3])) + 16'(A[0][2] * B[2][3])) + 16'(A[0][3] * B[3][3]);
    XOUT_[1][0] = (((0 + 16'(A[1][0] * B[0][0])) + 16'(A[1][1] * B[1][0])) + 16'(A[1][2] * B[2][0])) + 16'(A[1][3] * B[3][0]);
    XOUT_[1][1] = (((0 + 16'(A[1][0] * B[0][1])) + 16'(A[1][1] * B[1][1])) + 16'(A[1][2] * B[2][1])) + 16'(A[1][3] * B[3][1]);
    XOUT_[1][2] = (((0 + 16'(A[1][0] * B[0][2])) + 16'(A[1][1] * B[1][2])) + 16'(A[1][2] * B[2][2])) + 16'(A[1][3] * B[3][2]);
    XOUT_[1][3] = (((0 + 16'(A[1][0] * B[0][3])) + 16'(A[1][1] * B[1][3])) + 16'(A[1][2] * B[2][3])) + 16'(A[1][3] * B[3][3]);
    XOUT_[2][0] = (((0 + 16'(A[2][0] * B[0][0])) + 16'(A[2][1] * B[1][0])) + 16'(A[2][2] * B[2][0])) + 16'(A[2][3] * B[3][0]);
    XOUT_[2][1] = (((0 + 16'(A[2][0] * B[0][1])) + 16'(A[2][1] * B[1][1])) + 16'(A[2][2] * B[2][1])) + 16'(A[2][3] * B[3][1]);
    XOUT_[2][2] = (((0 + 16'(A[2][0] * B[0][2])) + 16'(A[2][1] * B[1][2])) + 16'(A[2][2] * B[2][2])) + 16'(A[2][3] * B[3][2]);
    XOUT_[2][3] = (((0 + 16'(A[2][0] * B[0][3])) + 16'(A[2][1] * B[1][3])) + 16'(A[2][2] * B[2][3])) + 16'(A[2][3] * B[3][3]);
    XOUT_[3][0] = (((0 + 16'(A[3][0] * B[0][0])) + 16'(A[3][1] * B[1][0])) + 16'(A[3][2] * B[2][0])) + 16'(A[3][3] * B[3][0]);
    XOUT_[3][1] = (((0 + 16'(A[3][0] * B[0][1])) + 16'(A[3][1] * B[1][1])) + 16'(A[3][2] * B[2][1])) + 16'(A[3][3] * B[3][1]);
    XOUT_[3][2] = (((0 + 16'(A[3][0] * B[0][2])) + 16'(A[3][1] * B[1][2])) + 16'(A[3][2] * B[2][2])) + 16'(A[3][3] * B[3][2]);
    XOUT_[3][3] = (((0 + 16'(A[3][0] * B[0][3])) + 16'(A[3][1] * B[1][3])) + 16'(A[3][2] * B[2][3])) + 16'(A[3][3] * B[3][3]);
  end
  assign XOUT = XOUT_;
endmodule
